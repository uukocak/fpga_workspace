library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity spi_ams is
    Port (
    CLK  : in  std_logic;
    LADC : out std_logic;
    SYNC : out std_logic;
    SCLK : out std_logic;
    DIN  : out std_logic
   -- out_test : out std_logic_vector(15 downto 0)
    );
end spi_ams;

architecture Behavioral of spi_ams is

    type state_t is (initialize, send_pack32, iterate_wave);
    type vector_array_t is array(0 to 359) of std_logic_vector(15 downto 0);

    signal state : state_t := initialize;
    signal package32 : std_logic_vector(31 downto 0);
    signal wave_array :  vector_array_t  :=  ( "1000000000000000",
    "1000001000111011",
    "1000010001110111",
    "1000011010110010",
    "1000100011101101",
    "1000101100100111",
    "1000110101100001",
    "1000111110011001",
    "1001000111010000",
    "1001010000000101",
    "1001011000111010",
    "1001100001101100",
    "1001101010011100",
    "1001110011001011",
    "1001111011110111",
    "1010000100100000",
    "1010001101000111",
    "1010010101101100",
    "1010011110001101",
    "1010100110101100",
    "1010101111000111",
    "1010110111011110",
    "1010111111110010",
    "1011001000000011",
    "1011010000001111",
    "1011011000011000",
    "1011100000011100",
    "1011101000011100",
    "1011110000010111",
    "1011111000001101",
    "1011111111111111",
    "1100000111101100",
    "1100001111010100",
    "1100010110110110",
    "1100011110010011",
    "1100100101101010",
    "1100101100111100",
    "1100110100000111",
    "1100111011001101",
    "1101000010001101",
    "1101001001000110",
    "1101001111111001",
    "1101010110100101",
    "1101011101001011",
    "1101100011101010",
    "1101101010000010",
    "1101110000010010",
    "1101110110011100",
    "1101111100011110",
    "1110000010011001",
    "1110001000001101",
    "1110001101111001",
    "1110010011011101",
    "1110011000111001",
    "1110011110001101",
    "1110100011011001",
    "1110101000011101",
    "1110101101011001",
    "1110110010001100",
    "1110110110110111",
    "1110111011011001",
    "1110111111110011",
    "1111000100000011",
    "1111001000001100",
    "1111001100001011",
    "1111010000000001",
    "1111010011101110",
    "1111010111010010",
    "1111011010101101",
    "1111011101111111",
    "1111100001000111",
    "1111100100000110",
    "1111100110111011",
    "1111101001100111",
    "1111101100001010",
    "1111101110100010",
    "1111110000110010",
    "1111110010110111",
    "1111110100110011",
    "1111110110100101",
    "1111111000001101",
    "1111111001101100",
    "1111111011000000",
    "1111111100001011",
    "1111111101001011",
    "1111111110000010",
    "1111111110101111",
    "1111111111010010",
    "1111111111101011",
    "1111111111111010",
    "1111111111111111",
    "1111111111111010",
    "1111111111101011",
    "1111111111010010",
    "1111111110101111",
    "1111111110000010",
    "1111111101001011",
    "1111111100001011",
    "1111111011000000",
    "1111111001101100",
    "1111111000001101",
    "1111110110100101",
    "1111110100110011",
    "1111110010110111",
    "1111110000110010",
    "1111101110100010",
    "1111101100001010",
    "1111101001100111",
    "1111100110111011",
    "1111100100000110",
    "1111100001000111",
    "1111011101111111",
    "1111011010101101",
    "1111010111010010",
    "1111010011101110",
    "1111010000000001",
    "1111001100001011",
    "1111001000001100",
    "1111000100000011",
    "1110111111110011",
    "1110111011011001",
    "1110110110110111",
    "1110110010001100",
    "1110101101011001",
    "1110101000011101",
    "1110100011011001",
    "1110011110001101",
    "1110011000111001",
    "1110010011011101",
    "1110001101111001",
    "1110001000001101",
    "1110000010011001",
    "1101111100011110",
    "1101110110011100",
    "1101110000010010",
    "1101101010000010",
    "1101100011101010",
    "1101011101001011",
    "1101010110100101",
    "1101001111111001",
    "1101001001000110",
    "1101000010001101",
    "1100111011001101",
    "1100110100000111",
    "1100101100111100",
    "1100100101101010",
    "1100011110010011",
    "1100010110110110",
    "1100001111010100",
    "1100000111101100",
    "1011111111111111",
    "1011111000001101",
    "1011110000010111",
    "1011101000011100",
    "1011100000011100",
    "1011011000011000",
    "1011010000001111",
    "1011001000000011",
    "1010111111110010",
    "1010110111011110",
    "1010101111000111",
    "1010100110101100",
    "1010011110001101",
    "1010010101101100",
    "1010001101000111",
    "1010000100100000",
    "1001111011110111",
    "1001110011001011",
    "1001101010011100",
    "1001100001101100",
    "1001011000111010",
    "1001010000000101",
    "1001000111010000",
    "1000111110011001",
    "1000110101100001",
    "1000101100100111",
    "1000100011101101",
    "1000011010110010",
    "1000010001110111",
    "1000001000111011",
    "1000000000000000",
    "0111110111000100",
    "0111101110001000",
    "0111100101001101",
    "0111011100010010",
    "0111010011011000",
    "0111001010011110",
    "0111000001100110",
    "0110111000101111",
    "0110101111111010",
    "0110100111000101",
    "0110011110010011",
    "0110010101100011",
    "0110001100110100",
    "0110000100001000",
    "0101111011011111",
    "0101110010111000",
    "0101101010010011",
    "0101100001110010",
    "0101011001010011",
    "0101010000111000",
    "0101001000100001",
    "0101000000001101",
    "0100110111111100",
    "0100101111110000",
    "0100100111100111",
    "0100011111100011",
    "0100010111100011",
    "0100001111101000",
    "0100000111110010",
    "0100000000000000",
    "0011111000010011",
    "0011110000101011",
    "0011101001001001",
    "0011100001101100",
    "0011011010010101",
    "0011010011000011",
    "0011001011111000",
    "0011000100110010",
    "0010111101110010",
    "0010110110111001",
    "0010110000000110",
    "0010101001011010",
    "0010100010110100",
    "0010011100010101",
    "0010010101111101",
    "0010001111101101",
    "0010001001100011",
    "0010000011100001",
    "0001111101100110",
    "0001110111110010",
    "0001110010000110",
    "0001101100100010",
    "0001100111000110",
    "0001100001110010",
    "0001011100100110",
    "0001010111100010",
    "0001010010100110",
    "0001001101110011",
    "0001001001001000",
    "0001000100100110",
    "0001000000001100",
    "0000111011111100",
    "0000110111110011",
    "0000110011110100",
    "0000101111111110",
    "0000101100010001",
    "0000101000101101",
    "0000100101010010",
    "0000100010000000",
    "0000011110111000",
    "0000011011111001",
    "0000011001000100",
    "0000010110011000",
    "0000010011110101",
    "0000010001011101",
    "0000001111001101",
    "0000001101001000",
    "0000001011001100",
    "0000001001011010",
    "0000000111110010",
    "0000000110010011",
    "0000000100111111",
    "0000000011110100",
    "0000000010110100",
    "0000000001111101",
    "0000000001010000",
    "0000000000101101",
    "0000000000010100",
    "0000000000000101",
    "0000000000000000",
    "0000000000000101",
    "0000000000010100",
    "0000000000101101",
    "0000000001010000",
    "0000000001111101",
    "0000000010110100",
    "0000000011110100",
    "0000000100111111",
    "0000000110010011",
    "0000000111110010",
    "0000001001011010",
    "0000001011001100",
    "0000001101001000",
    "0000001111001101",
    "0000010001011101",
    "0000010011110101",
    "0000010110011000",
    "0000011001000100",
    "0000011011111001",
    "0000011110111000",
    "0000100010000000",
    "0000100101010010",
    "0000101000101101",
    "0000101100010001",
    "0000101111111110",
    "0000110011110100",
    "0000110111110011",
    "0000111011111100",
    "0001000000001100",
    "0001000100100110",
    "0001001001001000",
    "0001001101110011",
    "0001010010100110",
    "0001010111100010",
    "0001011100100110",
    "0001100001110010",
    "0001100111000110",
    "0001101100100010",
    "0001110010000110",
    "0001110111110010",
    "0001111101100110",
    "0010000011100001",
    "0010001001100011",
    "0010001111101101",
    "0010010101111101",
    "0010011100010101",
    "0010100010110100",
    "0010101001011010",
    "0010110000000110",
    "0010110110111001",
    "0010111101110010",
    "0011000100110010",
    "0011001011111000",
    "0011010011000011",
    "0011011010010101",
    "0011100001101100",
    "0011101001001001",
    "0011110000101011",
    "0011111000010011",
    "0100000000000000",
    "0100000111110010",
    "0100001111101000",
    "0100010111100011",
    "0100011111100011",
    "0100100111100111",
    "0100101111110000",
    "0100110111111100",
    "0101000000001101",
    "0101001000100001",
    "0101010000111000",
    "0101011001010011",
    "0101100001110010",
    "0101101010010011",
    "0101110010111000",
    "0101111011011111",
    "0110000100001000",
    "0110001100110100",
    "0110010101100011",
    "0110011110010011",
    "0110100111000101",
    "0110101111111010",
    "0110111000101111",
    "0111000001100110",
    "0111001010011110",
    "0111010011011000",
    "0111011100010010",
    "0111100101001101",
    "0111101110001000",
    "0111110111000100"
);


    constant command : std_logic_vector(3 downto 0) := "0010";
    constant ch_addr : std_logic_vector(3 downto 0) := "0000";
    constant period : integer := 100; --nanoseconds

begin

    SCLK <= CLK;
    LADC <= '0';

    FSM : process(state,CLK)
        variable clk_counter : integer := 0;
        variable array_index : integer := 0;
        variable freq_coef : integer := 1;
    begin

        if ( CLK'event AND CLK = '1' ) then

            case(state) is

                when initialize =>
                    SYNC      <='1';
                    clk_counter := 0;
                    array_index := 0;
                    freq_coef   := 7;
                    state <= iterate_wave;

                when iterate_wave =>

                    if (clk_counter < 2000/period) then --Wait for 2us
                        state <= iterate_wave;
                        clk_counter := clk_counter + 1;
                    else
                        if(array_index > 359) then
                            array_index := array_index-360;
                            package32 <= "0000" & command & ch_addr & wave_array(array_index) & "0000";
                        else
                            package32 <= "0000" & command & ch_addr & wave_array(array_index) & "0000";
                        end if;
                        clk_counter := clk_counter + 1;
                        --out_test <= wave_array(array_index); --test
                        array_index := array_index + freq_coef;
                        state <= send_pack32;
                        clk_counter := 0;
                    end if;


                when send_pack32 =>
                    if ( clk_counter < 32 ) then
                        SYNC <= '0';
                        DIN    <= package32(31-clk_counter);
                        state  <= send_pack32;
                        clk_counter := clk_counter + 1;
                    else
                        SYNC <= '1';
                        DIN    <= '0';
                        state  <= iterate_wave;
                        clk_counter := 0;
                    end if;


                when others =>

            end case;

        end if;


    end process;


end Behavioral;
