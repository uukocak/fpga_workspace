library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity spi_ams is
    Port (
    CLK  : in  std_logic;
    LADC : out std_logic;
    SYNC : out std_logic;
    SCLK : out std_logic;
    DIN  : out std_logic
   -- out_test : out std_logic_vector(15 downto 0)
    );
end spi_ams;

architecture Behavioral of spi_ams is

    type state_t is (initialize, send_pack32, iterate_wave);
    type vector_array_t is array(0 to 359) of std_logic_vector(15 downto 0);

    signal state : state_t := initialize;
    signal package32 : std_logic_vector(31 downto 0);
    signal wave_array :  vector_array_t  :=  ( "011001100110011",
    "011010000011000",
    "011010011111100",
    "011010111100001",
    "011011011000101",
    "011011110101001",
    "011100010001101",
    "011100101110000",
    "011101001010011",
    "011101100110101",
    "011110000010111",
    "011110011111000",
    "011110111011000",
    "011111010110111",
    "011111110010110",
    "100000001110011",
    "100000101010000",
    "100001000101011",
    "100001100000101",
    "100001111011110",
    "100010010110110",
    "100010110001100",
    "100011001100001",
    "100011100110100",
    "100100000000110",
    "100100011010110",
    "100100110100101",
    "100101001110001",
    "100101100111100",
    "100110000000101",
    "100110011001100",
    "100110110010010",
    "100111001010101",
    "100111100010110",
    "100111111010100",
    "101000010010001",
    "101000101001011",
    "101001000000011",
    "101001010111000",
    "101001101101100",
    "101010000011100",
    "101010011001010",
    "101010101110101",
    "101011000011110",
    "101011011000100",
    "101011101100111",
    "101100000000111",
    "101100010100101",
    "101100100111111",
    "101100111010111",
    "101101001101100",
    "101101011111101",
    "101101110001011",
    "101110000010111",
    "101110010011111",
    "101110100100100",
    "101110110100101",
    "101111000100011",
    "101111010011110",
    "101111100010110",
    "101111110001010",
    "101111111111011",
    "110000001101000",
    "110000011010001",
    "110000100110111",
    "110000110011010",
    "110000111111001",
    "110001001010100",
    "110001010101100",
    "110001011111111",
    "110001101010000",
    "110001110011100",
    "110001111100100",
    "110010000101001",
    "110010001101010",
    "110010010100111",
    "110010011100001",
    "110010100010110",
    "110010101001000",
    "110010101110101",
    "110010110011111",
    "110010111000101",
    "110010111100110",
    "110011000000100",
    "110011000011110",
    "110011000110100",
    "110011001000110",
    "110011001010100",
    "110011001011110",
    "110011001100100",
    "110011001100110",
    "110011001100100",
    "110011001011110",
    "110011001010100",
    "110011001000110",
    "110011000110100",
    "110011000011110",
    "110011000000100",
    "110010111100110",
    "110010111000101",
    "110010110011111",
    "110010101110101",
    "110010101001000",
    "110010100010110",
    "110010011100001",
    "110010010100111",
    "110010001101010",
    "110010000101001",
    "110001111100100",
    "110001110011100",
    "110001101010000",
    "110001011111111",
    "110001010101100",
    "110001001010100",
    "110000111111001",
    "110000110011010",
    "110000100110111",
    "110000011010001",
    "110000001101000",
    "101111111111011",
    "101111110001010",
    "101111100010110",
    "101111010011110",
    "101111000100011",
    "101110110100101",
    "101110100100100",
    "101110010011111",
    "101110000010111",
    "101101110001011",
    "101101011111101",
    "101101001101100",
    "101100111010111",
    "101100100111111",
    "101100010100101",
    "101100000000111",
    "101011101100111",
    "101011011000100",
    "101011000011110",
    "101010101110101",
    "101010011001010",
    "101010000011100",
    "101001101101100",
    "101001010111000",
    "101001000000011",
    "101000101001011",
    "101000010010001",
    "100111111010100",
    "100111100010110",
    "100111001010101",
    "100110110010010",
    "100110011001101",
    "100110000000101",
    "100101100111100",
    "100101001110001",
    "100100110100101",
    "100100011010110",
    "100100000000110",
    "100011100110100",
    "100011001100001",
    "100010110001100",
    "100010010110110",
    "100001111011110",
    "100001100000101",
    "100001000101011",
    "100000101010000",
    "100000001110011",
    "011111110010110",
    "011111010110111",
    "011110111011000",
    "011110011111000",
    "011110000010111",
    "011101100110101",
    "011101001010011",
    "011100101110000",
    "011100010001101",
    "011011110101001",
    "011011011000101",
    "011010111100001",
    "011010011111100",
    "011010000011000",
    "011001100110011",
    "011001001001110",
    "011000101101010",
    "011000010000101",
    "010111110100001",
    "010111010111101",
    "010110111011001",
    "010110011110110",
    "010110000010011",
    "010101100110001",
    "010101001001111",
    "010100101101110",
    "010100010001110",
    "010011110101111",
    "010011011010000",
    "010010111110011",
    "010010100010110",
    "010010000111011",
    "010001101100001",
    "010001010001000",
    "010000110110000",
    "010000011011010",
    "010000000000101",
    "001111100110010",
    "001111001100000",
    "001110110010000",
    "001110011000001",
    "001101111110101",
    "001101100101010",
    "001101001100001",
    "001100110011010",
    "001100011010100",
    "001100000010001",
    "001011101010000",
    "001011010010010",
    "001010111010101",
    "001010100011011",
    "001010001100011",
    "001001110101110",
    "001001011111010",
    "001001001001010",
    "001000110011100",
    "001000011110001",
    "001000001001000",
    "000111110100010",
    "000111011111111",
    "000111001011111",
    "000110111000001",
    "000110100100111",
    "000110010001111",
    "000101111111010",
    "000101101101001",
    "000101011011011",
    "000101001001111",
    "000100111000111",
    "000100101000010",
    "000100011000001",
    "000100001000011",
    "000011111001000",
    "000011101010000",
    "000011011011100",
    "000011001101011",
    "000010111111110",
    "000010110010101",
    "000010100101111",
    "000010011001100",
    "000010001101101",
    "000010000010010",
    "000001110111010",
    "000001101100111",
    "000001100010110",
    "000001011001010",
    "000001010000010",
    "000001000111101",
    "000000111111100",
    "000000110111111",
    "000000110000101",
    "000000101010000",
    "000000100011110",
    "000000011110001",
    "000000011000111",
    "000000010100001",
    "000000010000000",
    "000000001100010",
    "000000001001000",
    "000000000110010",
    "000000000100000",
    "000000000010010",
    "000000000001000",
    "000000000000010",
    "000000000000000",
    "000000000000010",
    "000000000001000",
    "000000000010010",
    "000000000100000",
    "000000000110010",
    "000000001001000",
    "000000001100010",
    "000000010000000",
    "000000010100001",
    "000000011000111",
    "000000011110001",
    "000000100011110",
    "000000101010000",
    "000000110000101",
    "000000110111111",
    "000000111111100",
    "000001000111101",
    "000001010000010",
    "000001011001010",
    "000001100010110",
    "000001101100111",
    "000001110111010",
    "000010000010010",
    "000010001101101",
    "000010011001100",
    "000010100101111",
    "000010110010101",
    "000010111111110",
    "000011001101011",
    "000011011011100",
    "000011101010000",
    "000011111001000",
    "000100001000011",
    "000100011000001",
    "000100101000010",
    "000100111000111",
    "000101001001111",
    "000101011011011",
    "000101101101001",
    "000101111111010",
    "000110010001111",
    "000110100100111",
    "000110111000001",
    "000111001011111",
    "000111011111111",
    "000111110100010",
    "001000001001000",
    "001000011110001",
    "001000110011100",
    "001001001001010",
    "001001011111010",
    "001001110101110",
    "001010001100011",
    "001010100011011",
    "001010111010101",
    "001011010010010",
    "001011101010000",
    "001100000010001",
    "001100011010100",
    "001100110011001",
    "001101001100001",
    "001101100101010",
    "001101111110101",
    "001110011000001",
    "001110110010000",
    "001111001100000",
    "001111100110010",
    "010000000000101",
    "010000011011010",
    "010000110110000",
    "010001010001000",
    "010001101100001",
    "010010000111011",
    "010010100010110",
    "010010111110011",
    "010011011010000",
    "010011110101111",
    "010100010001110",
    "010100101101110",
    "010101001001111",
    "010101100110001",
    "010110000010011",
    "010110011110110",
    "010110111011001",
    "010111010111101",
    "010111110100001",
    "011000010000101",
    "011000101101010",
    "011001001001110"
);

    constant command : std_logic_vector(3 downto 0) := "0010";
    constant ch_addr : std_logic_vector(3 downto 0) := "0011";
    constant period : integer := 200; --nanoseconds

begin

    SCLK <= CLK;
    LADC <= '0';

    FSM : process(state,CLK)
        variable clk_counter : integer := 0;
        variable array_index : integer := 0;
        variable freq_coef : integer := 1;
    begin

        if ( CLK'event AND CLK = '1' ) then

            case(state) is

                when initialize =>
                    SYNC      <='1';
                    clk_counter := 0;
                    array_index := 0;
                    freq_coef   := 1;
                    state <= iterate_wave;

                when iterate_wave =>

                    if (clk_counter < 100000/period) then --Wait for 2us
                        state <= iterate_wave;
                        clk_counter := clk_counter + 1;
                    else
                        if(array_index > 359) then
                            array_index := array_index-360;
                            package32 <= "0000" & command & ch_addr & wave_array(array_index) & "0000";
                        else
                            package32 <= "0000" & command & ch_addr & wave_array(array_index) & "0000";
                        end if;
                        --out_test <= wave_array(array_index); --test
                        array_index := array_index + freq_coef;
                        state <= send_pack32;
                        clk_counter := 0;
                    end if;


                when send_pack32 =>
                    if ( clk_counter < 32 ) then
                        SYNC <= '0';
                        DIN    <= package32(31-clk_counter);
                        state  <= send_pack32;
                        clk_counter := clk_counter + 1;
                    else
                        SYNC <= '1';
                        DIN    <= '0';
                        state  <= iterate_wave;
                        clk_counter := 0;
                    end if;


                when others =>

            end case;

        end if;


    end process;


end Behavioral;
